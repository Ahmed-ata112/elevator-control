-- 2 modules should exist in here 